`timescale 1ns / 1ps


module filter #(parameter NR_STAGES = 32,
				parameter DWIDTH = 16,
				parameter DDWIDTH = 2*DWIDTH,
				parameter CWIDTH = NR_STAGES * DWIDTH)
			   (input  clk,
				input  rst,
				output req_in,
				input  ack_in,
				input  [0:DWIDTH-1] data_in,
				output req_out,
				input  ack_out,
				output [0:DWIDTH-1] data_out,
				input  [0:CWIDTH-1] h_in);

	// Output request register
	reg req_out_buf;
	assign req_out = req_out_buf;

	// Input request register
	reg req_in_buf;
	assign req_in = req_in_buf;
  
	reg [0:5] stage; // Counter for the stage we're in
	reg signed [0:DWIDTH-1] in [0:NR_STAGES-1]; // Cached inputs
	reg signed [0:DDWIDTH-1] sum; // Accumulator
	reg signed [0:DDWIDTH-1] acc; // Accumulator
	reg signed [0:DWIDTH-1] out;
	assign data_out = out;

	reg [0:5] i;

	always @(posedge clk)
	begin
		// Reset => initialize
		if (rst)
		begin
			req_in_buf <= 0;
			req_out_buf <= 0;
			sum <= 0;
			acc <= 0;
			stage <= 0;
		end
		// !Reset => run
		else
		begin
			// Input request & acknowledge => read input and signal input done
			if (req_in && ack_in)
			begin
				sum <= 0;
				acc <= 0;
				in[0] <= data_in;
				for (i = 0; i < NR_STAGES - 1; i = i + 1)
				begin
					in[i + 1] <= in[i];
				end
				req_in_buf <= 0;
			end
			// Output request & acknowledge => signal output done
			if (req_out && ack_out)
			begin
				req_out_buf <= 0;
			end
			// If we need no inputs and have no outputs ready, and are out of startup phase
			// then proceed with the computation
			if (!req_in && !req_out && !ack_in && !ack_out)
			begin   
				if (stage == NR_STAGES)
				begin
					req_in_buf <= 1;
					req_out_buf <= 1;
					out <= sum + acc;
					stage <= 0;
				end
				else
				begin
					acc <= (in[stage] * $signed(h_in[stage*DWIDTH+:DWIDTH])) >> DWIDTH;
					sum <= sum + acc;
					stage <= stage + 1;
				end
			end
		end
	end

endmodule
